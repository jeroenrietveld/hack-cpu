-------------------------------------------------------------------------------
-- Title      : Testbench for design "alu"
-- Project    :
-------------------------------------------------------------------------------
-- File       : alu_tb.vhd
-- Author     : Jeroen Rietveld  <jeroenrietveld@Macbook-Pro-Jeroen.local>
-- Company    :
-- Created    : 2019-07-08
-- Last update: 2019-07-09
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------
-- Copyright (c) 2019
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-07-08  1.0      jeroenrietveld  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------------

entity alu_tb is

end entity alu_tb;

-------------------------------------------------------------------------------

architecture arch of alu_tb is

  -- component ports
  signal I_A          : std_logic_vector(15 downto 0);
  signal I_B          : std_logic_vector(15 downto 0);
  signal I_zeroA      : std_logic;
  signal I_zeroB      : std_logic;
  signal I_notA       : std_logic;
  signal I_notB       : std_logic;
  signal I_function   : std_logic;
  signal I_notO       : std_logic;
  signal O_out        : std_logic_vector(15 downto 0);
  signal O_zero       : std_logic;
  signal O_notGreater : std_logic;

  -- clock
  signal Clk          : std_logic := '1';
  constant clk_period : time      := 20 ns;
begin  -- architecture arch

  -- component instantiation
  DUT : entity work.alu
    port map (
      I_A          => I_A,
      I_B          => I_B,
      I_zeroA      => I_zeroA,
      I_zeroB      => I_zeroB,
      I_notA       => I_notA,
      I_notB       => I_notB,
      I_function   => I_function,
      I_notO       => I_notO,
      O_out        => O_out,
      O_zero       => O_zero,
      O_notGreater => O_notGreater);

  -- clock generation
  Clk <= not Clk after 10 ns;
  process
    type pattern_type is record
      --  The inputs of the alu.
      x, y                  : std_logic_vector(15 downto 0);
      zx, nx, zy, ny, f, no : std_logic;
      --  The expected outputs of the alu.
      cout                  : std_logic_vector(15 downto 0);
      zr, ng                : std_logic;
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array :=
        (("0000000000000000", "1111111111111111", '1', '0', '1', '0', '1', '0', "0000000000000000", '1', '0'),
         ("0000000000000000", "1111111111111111", '1', '1', '1', '1', '1', '1', "0000000000000001", '0', '0'),
         ("0000000000000000", "1111111111111111", '1', '1', '1', '0', '1', '0', "1111111111111111", '0', '1'),
         ("0000000000000000", "1111111111111111", '0', '0', '1', '1', '0', '0', "0000000000000000", '1', '0'),
         ("0000000000000000", "1111111111111111", '1', '1', '0', '0', '0', '0', "1111111111111111", '0', '1'),
         ("0000000000000000", "1111111111111111", '0', '0', '1', '1', '0', '1', "1111111111111111", '0', '1'),
         ("0000000000000000", "1111111111111111", '1', '1', '0', '0', '0', '1', "0000000000000000", '1', '0'),
         ("0000000000000000", "1111111111111111", '0', '0', '1', '1', '1', '1', "0000000000000000", '1', '0'),
         ("0000000000000000", "1111111111111111", '1', '1', '0', '0', '1', '1', "0000000000000001", '0', '0'),
         ("0000000000000000", "1111111111111111", '0', '1', '1', '1', '1', '1', "0000000000000001", '0', '0'),
         ("0000000000000000", "1111111111111111", '1', '1', '0', '1', '1', '1', "0000000000000000", '1', '0'),
         ("0000000000000000", "1111111111111111", '0', '0', '1', '1', '1', '0', "1111111111111111", '0', '1'),
         ("0000000000000000", "1111111111111111", '1', '1', '0', '0', '1', '0', "1111111111111110", '0', '1'),
         ("0000000000000000", "1111111111111111", '0', '0', '0', '0', '1', '0', "1111111111111111", '0', '1'),
         ("0000000000000000", "1111111111111111", '0', '1', '0', '0', '1', '1', "0000000000000001", '0', '0'),
         ("0000000000000000", "1111111111111111", '0', '0', '0', '1', '1', '1', "1111111111111111", '0', '1'),
         ("0000000000000000", "1111111111111111", '0', '0', '0', '0', '0', '0', "0000000000000000", '1', '0'),
         ("0000000000000000", "1111111111111111", '0', '1', '0', '1', '0', '1', "1111111111111111", '0', '1'),
         ("0000000000010001", "0000000000000011", '1', '0', '1', '0', '1', '0', "0000000000000000", '1', '0'),
         ("0000000000010001", "0000000000000011", '1', '1', '1', '1', '1', '1', "0000000000000001", '0', '0'),
         ("0000000000010001", "0000000000000011", '1', '1', '1', '0', '1', '0', "1111111111111111", '0', '1'),
         ("0000000000010001", "0000000000000011", '0', '0', '1', '1', '0', '0', "0000000000010001", '0', '0'),
         ("0000000000010001", "0000000000000011", '1', '1', '0', '0', '0', '0', "0000000000000011", '0', '0'),
         ("0000000000010001", "0000000000000011", '0', '0', '1', '1', '0', '1', "1111111111101110", '0', '1'),
         ("0000000000010001", "0000000000000011", '1', '1', '0', '0', '0', '1', "1111111111111100", '0', '1'),
         ("0000000000010001", "0000000000000011", '0', '0', '1', '1', '1', '1', "1111111111101111", '0', '1'),
         ("0000000000010001", "0000000000000011", '1', '1', '0', '0', '1', '1', "1111111111111101", '0', '1'),
         ("0000000000010001", "0000000000000011", '0', '1', '1', '1', '1', '1', "0000000000010010", '0', '0'),
         ("0000000000010001", "0000000000000011", '1', '1', '0', '1', '1', '1', "0000000000000100", '0', '0'),
         ("0000000000010001", "0000000000000011", '0', '0', '1', '1', '1', '0', "0000000000010000", '0', '0'),
         ("0000000000010001", "0000000000000011", '1', '1', '0', '0', '1', '0', "0000000000000010", '0', '0'),
         ("0000000000010001", "0000000000000011", '0', '0', '0', '0', '1', '0', "0000000000010100", '0', '0'),
         ("0000000000010001", "0000000000000011", '0', '1', '0', '0', '1', '1', "0000000000001110", '0', '0'),
         ("0000000000010001", "0000000000000011", '0', '0', '0', '1', '1', '1', "1111111111110010", '0', '1'),
         ("0000000000010001", "0000000000000011", '0', '0', '0', '0', '0', '0', "0000000000000001", '0', '0'),
         ("0000000000010001", "0000000000000011", '0', '1', '0', '1', '0', '1', "0000000000010011", '0', '0'));
  begin
    wait for clk_period;
    wait for clk_period/2;

    for i in patterns'range loop
      --  Set the inputs.
      I_A        <= patterns(i).x;
      I_B        <= patterns(i).y;
      I_zeroA    <= patterns(i).zx;
      I_notA     <= patterns(i).nx;
      I_zeroB    <= patterns(i).zy;
      I_notB     <= patterns(i).ny;
      I_function <= patterns(i).f;
      I_notO     <= patterns(i).no;

      wait for 1 ns;

      assert O_out = patterns(i).cout
        report "Incorrect O_data, expected " & integer'image(to_integer(signed(patterns(i).cout))) &
        " but got " & integer'image(to_integer(signed(O_out))) &
        " on iteration " & integer'image(i)
        severity error;

      -- assert O_zero = patterns(i).zr
      --   report "Incorrect O_data, expected " & integer'image(to_integer(signed(patterns(i).cout))) &
      --   " but got " & integer'image(to_integer(signed(O_zero)))
      --   severity error;

      -- assert O_notGreater = patterns(i).ng
      --   report "Incorrect O_data, expected " & integer'image(to_integer(signed(patterns(i).ng))) &
      --   " but got " & integer'image(to_integer(signed(O_notGreater)))
      --   severity error;

      wait for clk_period - 1 ns;
    end loop;

    assert false report "end of test" severity failure;
  end process;
end architecture arch;

-------------------------------------------------------------------------------

-- configuration alu_tb_arch_cfg of alu_tb is
-- end alu_tb_arch_cfg;

-------------------------------------------------------------------------------
