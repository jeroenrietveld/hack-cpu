-------------------------------------------------------------------------------
-- Title      : Testbench for design "ram16_n"
-- Project    :
-------------------------------------------------------------------------------
-- File       : ram16_n_tb.vhd
-- Author     : Jeroen Rietveld  <jeroenrietveld@Macbook-Pro-Jeroen.local>
-- Company    :
-- Created    : 2019-07-05
-- Last update: 2019-07-05
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------
-- Copyright (c) 2019
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-07-05  1.0      jeroenrietveld  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------------

entity ram16_n_tb is

end entity ram16_n_tb;

-------------------------------------------------------------------------------

architecture arch of ram16_n_tb is

  -- component generics
  constant N : positive := 8;

  -- component ports
  signal I_clk  : std_logic;
  signal I_data : std_logic_vector(15 downto 0);
  signal I_addr : natural;
  signal I_load : std_logic;
  signal O_data : std_logic_vector(15 downto 0);

  -- clock
  signal Clk          : std_logic := '1';
  constant clk_period : time      := 20 ns;
begin  -- architecture arch

  -- component instantiation
  DUT : entity work.ram16_n
    generic map (
      N => N)
    port map (
      I_clk  => Clk,
      I_data => I_data,
      I_addr => I_addr,
      I_load => I_load,
      O_data => O_data);

  -- clock generation
  Clk <= not Clk after clk_period / 2;

  process
    type pattern_type is record
      I_data : std_logic_vector(15 downto 0);
      I_load : std_logic;
      I_addr : std_logic_vector(2 downto 0);
      --  The output of the ram8.
      O_data : std_logic_vector(15 downto 0);
      -- I_data, I_addr : integer;
      -- I_load         : std_logic;
      -- O_data         : integer;
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array :=
              (("0000000000000000", '0', "000", "0000000000000000"),
         ("0000000000000000", '0', "000", "0000000000000000"),
         ("0000000000000000", '1', "000", "0000000000000000"),
         ("0000000000000000", '1', "000", "0000000000000000"),
         ("0010101101100111", '0', "000", "0000000000000000"),
         ("0010101101100111", '0', "000", "0000000000000000"),
         ("0010101101100111", '1', "001", "0000000000000000"),
         ("0010101101100111", '1', "001", "0010101101100111"),
         ("0010101101100111", '0', "000", "0000000000000000"),
         ("0010101101100111", '0', "000", "0000000000000000"),
         ("0000110100000101", '0', "011", "0000000000000000"),
         ("0000110100000101", '0', "011", "0000000000000000"),
         ("0000110100000101", '1', "011", "0000000000000000"),
         ("0000110100000101", '1', "011", "0000110100000101"),
         ("0000110100000101", '0', "011", "0000110100000101"),
         ("0000110100000101", '0', "011", "0000110100000101"),
         ("0000110100000101", '0', "001", "0010101101100111"),
         ("0001111001100001", '0', "001", "0010101101100111"),
         ("0001111001100001", '0', "001", "0010101101100111"),
         ("0001111001100001", '1', "111", "0000000000000000"),
         ("0001111001100001", '1', "111", "0001111001100001"),
         ("0001111001100001", '0', "111", "0001111001100001"),
         ("0001111001100001", '0', "111", "0001111001100001"),
         ("0001111001100001", '0', "011", "0000110100000101"),
         ("0001111001100001", '0', "111", "0001111001100001"),
         ("0001111001100001", '0', "000", "0000000000000000"),
         ("0001111001100001", '0', "000", "0000000000000000"),
         ("0001111001100001", '0', "001", "0010101101100111"),
         ("0001111001100001", '0', "010", "0000000000000000"),
         ("0001111001100001", '0', "011", "0000110100000101"),
         ("0001111001100001", '0', "100", "0000000000000000"),
         ("0001111001100001", '0', "101", "0000000000000000"),
         ("0001111001100001", '0', "110", "0000000000000000"),
         ("0001111001100001", '0', "111", "0001111001100001"),
         ("0101010101010101", '1', "000", "0000000000000000"),
         ("0101010101010101", '1', "000", "0101010101010101"),
         ("0101010101010101", '1', "001", "0010101101100111"),
         ("0101010101010101", '1', "001", "0101010101010101"),
         ("0101010101010101", '1', "010", "0000000000000000"),
         ("0101010101010101", '1', "010", "0101010101010101"),
         ("0101010101010101", '1', "011", "0000110100000101"),
         ("0101010101010101", '1', "011", "0101010101010101"),
         ("0101010101010101", '1', "100", "0000000000000000"),
         ("0101010101010101", '1', "100", "0101010101010101"),
         ("0101010101010101", '1', "101", "0000000000000000"),
         ("0101010101010101", '1', "101", "0101010101010101"),
         ("0101010101010101", '1', "110", "0000000000000000"),
         ("0101010101010101", '1', "110", "0101010101010101"),
         ("0101010101010101", '1', "111", "0001111001100001"),
         ("0101010101010101", '1', "111", "0101010101010101"),
         ("0101010101010101", '0', "000", "0101010101010101"),
         ("0101010101010101", '0', "000", "0101010101010101"),
         ("0101010101010101", '0', "001", "0101010101010101"),
         ("0101010101010101", '0', "010", "0101010101010101"),
         ("0101010101010101", '0', "011", "0101010101010101"),
         ("0101010101010101", '0', "100", "0101010101010101"),
         ("0101010101010101", '0', "101", "0101010101010101"),
         ("0101010101010101", '0', "110", "0101010101010101"),
         ("0101010101010101", '0', "111", "0101010101010101"),
         ("0101010101010110", '1', "000", "0101010101010101"),
         ("0101010101010110", '1', "000", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010110"),
         ("0101010101010110", '0', "001", "0101010101010101"),
         ("0101010101010110", '0', "010", "0101010101010101"),
         ("0101010101010110", '0', "011", "0101010101010101"),
         ("0101010101010110", '0', "100", "0101010101010101"),
         ("0101010101010110", '0', "101", "0101010101010101"),
         ("0101010101010110", '0', "110", "0101010101010101"),
         ("0101010101010110", '0', "111", "0101010101010101"),
         ("0101010101010101", '1', "000", "0101010101010110"),
         ("0101010101010101", '1', "000", "0101010101010101"),
         ("0101010101010110", '1', "001", "0101010101010101"),
         ("0101010101010110", '1', "001", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "001", "0101010101010110"),
         ("0101010101010110", '0', "010", "0101010101010101"),
         ("0101010101010110", '0', "011", "0101010101010101"),
         ("0101010101010110", '0', "100", "0101010101010101"),
         ("0101010101010110", '0', "101", "0101010101010101"),
         ("0101010101010110", '0', "110", "0101010101010101"),
         ("0101010101010110", '0', "111", "0101010101010101"),
         ("0101010101010101", '1', "001", "0101010101010110"),
         ("0101010101010101", '1', "001", "0101010101010101"),
         ("0101010101010110", '1', "010", "0101010101010101"),
         ("0101010101010110", '1', "010", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "001", "0101010101010101"),
         ("0101010101010110", '0', "010", "0101010101010110"),
         ("0101010101010110", '0', "011", "0101010101010101"),
         ("0101010101010110", '0', "100", "0101010101010101"),
         ("0101010101010110", '0', "101", "0101010101010101"),
         ("0101010101010110", '0', "110", "0101010101010101"),
         ("0101010101010110", '0', "111", "0101010101010101"),
         ("0101010101010101", '1', "010", "0101010101010110"),
         ("0101010101010101", '1', "010", "0101010101010101"),
         ("0101010101010110", '1', "011", "0101010101010101"),
         ("0101010101010110", '1', "011", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "001", "0101010101010101"),
         ("0101010101010110", '0', "010", "0101010101010101"),
         ("0101010101010110", '0', "011", "0101010101010110"),
         ("0101010101010110", '0', "100", "0101010101010101"),
         ("0101010101010110", '0', "101", "0101010101010101"),
         ("0101010101010110", '0', "110", "0101010101010101"),
         ("0101010101010110", '0', "111", "0101010101010101"),
         ("0101010101010101", '1', "011", "0101010101010110"),
         ("0101010101010101", '1', "011", "0101010101010101"),
         ("0101010101010110", '1', "100", "0101010101010101"),
         ("0101010101010110", '1', "100", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "001", "0101010101010101"),
         ("0101010101010110", '0', "010", "0101010101010101"),
         ("0101010101010110", '0', "011", "0101010101010101"),
         ("0101010101010110", '0', "100", "0101010101010110"),
         ("0101010101010110", '0', "101", "0101010101010101"),
         ("0101010101010110", '0', "110", "0101010101010101"),
         ("0101010101010110", '0', "111", "0101010101010101"),
         ("0101010101010101", '1', "100", "0101010101010110"),
         ("0101010101010101", '1', "100", "0101010101010101"),
         ("0101010101010110", '1', "101", "0101010101010101"),
         ("0101010101010110", '1', "101", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "001", "0101010101010101"),
         ("0101010101010110", '0', "010", "0101010101010101"),
         ("0101010101010110", '0', "011", "0101010101010101"),
         ("0101010101010110", '0', "100", "0101010101010101"),
         ("0101010101010110", '0', "101", "0101010101010110"),
         ("0101010101010110", '0', "110", "0101010101010101"),
         ("0101010101010110", '0', "111", "0101010101010101"),
         ("0101010101010101", '1', "101", "0101010101010110"),
         ("0101010101010101", '1', "101", "0101010101010101"),
         ("0101010101010110", '1', "110", "0101010101010101"),
         ("0101010101010110", '1', "110", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "001", "0101010101010101"),
         ("0101010101010110", '0', "010", "0101010101010101"),
         ("0101010101010110", '0', "011", "0101010101010101"),
         ("0101010101010110", '0', "100", "0101010101010101"),
         ("0101010101010110", '0', "101", "0101010101010101"),
         ("0101010101010110", '0', "110", "0101010101010110"),
         ("0101010101010110", '0', "111", "0101010101010101"),
         ("0101010101010101", '1', "110", "0101010101010110"),
         ("0101010101010101", '1', "110", "0101010101010101"),
         ("0101010101010110", '1', "111", "0101010101010101"),
         ("0101010101010110", '1', "111", "0101010101010110"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "000", "0101010101010101"),
         ("0101010101010110", '0', "001", "0101010101010101"),
         ("0101010101010110", '0', "010", "0101010101010101"),
         ("0101010101010110", '0', "011", "0101010101010101"),
         ("0101010101010110", '0', "100", "0101010101010101"),
         ("0101010101010110", '0', "101", "0101010101010101"),
         ("0101010101010110", '0', "110", "0101010101010101"),
         ("0101010101010110", '0', "111", "0101010101010110"),
         ("0101010101010101", '1', "111", "0101010101010110"),
         ("0101010101010101", '1', "111", "0101010101010101"),
         ("0101010101010101", '0', "000", "0101010101010101"),
         ("0101010101010101", '0', "000", "0101010101010101"),
         ("0101010101010101", '0', "001", "0101010101010101"),
         ("0101010101010101", '0', "010", "0101010101010101"),
         ("0101010101010101", '0', "011", "0101010101010101"),
         ("0101010101010101", '0', "100", "0101010101010101"),
         ("0101010101010101", '0', "101", "0101010101010101"),
         ("0101010101010101", '0', "110", "0101010101010101"),
         ("0101010101010101", '0', "111", "0101010101010101"));
  begin
    wait for clk_period;
    wait for clk_period/2;

    for i in patterns'range loop
      -- I_data <= std_logic_vector(to_signed(patterns(i).I_data, I_data'length));
      I_data <= patterns(i).I_data;
      I_addr <= to_integer(unsigned(patterns(i).I_addr));
      I_load <= patterns(i).I_load;

      wait for 1 ns;

      -- assert O_data = std_logic_vector(to_signed(patterns(i).O_data, O_data'length))
      assert O_data = patterns(i).O_data
        report "Incorrect O_data, expected " & integer'image(to_integer(signed(patterns(i).O_data))) &
        " but got " & integer'image(to_integer(signed(O_data))) &
        " for address " & integer'image(to_integer(unsigned(patterns(i).I_addr))) &
        " on iteration " & integer'image(i)
        severity error;

      wait for clk_period - 1 ns;
    end loop;

    assert false report "end of test" severity failure;
  end process;
end arch;

-------------------------------------------------------------------------------

configuration ram16_n_tb_arch_cfg of ram16_n_tb is
  for arch
  end for;
end ram16_n_tb_arch_cfg;

-------------------------------------------------------------------------------
